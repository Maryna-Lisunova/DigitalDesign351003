library ieee;
use ieee.std_logic_1164.all;

entity task7 is
    port (
    led_o: out std_logic_vector(15 downto 0);
    sw_i: in std_logic_vector(15 downto 0)
    );
end task7;

architecture rtl of task7 is
begin

end rtl;